library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.math_real.all;

library work;
use work.basic.all;
use work.add.all;

entity data_path is
  port (
    
  ) ;
end data_path;
--- Control Signals

-- Instruction Register
----- wr_enable


architecture flow of data_path is


begin


end flow;