library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all;
use ieee.numeric_std.all;

-- Package Declarations
package elem is
    component reg_ent is
        port(  );
    end component;
end package;

-- Entity and Architecture Declarations
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


